
module aes_top(
	input 
);
