module AddRoundKey(
	input [0:127] i_plain,
	input []
);