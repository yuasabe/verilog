module SubBytes(
	input 
);