module ShiftRows(
	input i_clock,
	input [0:127] i_data,
	input i_active,
	output [0:127] o_data
);

endmodule